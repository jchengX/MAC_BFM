package mac_pkg;
  import uvm_pkg::*;
  
  `include "mac_sequencer.sv"
  `include "mac_monitor.sv"
  `include "mac_driver.sv"
  `include "mac_agent.sv"
  `include "mac_scoreboard.sv"
  `include "mac_config.sv"
  `include "mac_env.sv"
  `include "mac_test.sv"
endpackage: mac_pkg
