class data_packet
