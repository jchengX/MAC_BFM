class beacon_packet extends packet;

  
