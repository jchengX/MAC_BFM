package crc7_pkg;
  import uvm_pkg::*;
  
  `include "crc7_sequencer.sv"
  `include "crc7_monitor.sv"
  `include "crc7_driver.sv"
  `include "crc7_agent.sv"
  `include "crc7_scoreboard.sv"
  `include "crc7_config.sv"
  `include "crc7_env.sv"
  `include "crc7_test.sv"
endpackage: crc7_pkg
