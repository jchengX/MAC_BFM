class aggregate_packet
