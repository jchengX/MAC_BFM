class beacon_packet extends packet;
  type = 2'b00;
  sub_type = 4'b1000;
  

  
